module DP_DDR3();

endmodule